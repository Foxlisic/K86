/**
 * Здесь исполняются инструкции
 */

always @(posedge clock)
begin

end
