`timescale 10ns / 1ns
module tb;
// -----------------------------------------------------------------------------
reg         clock, reset_n;
always #2.0 clock = ~clock;
// -----------------------------------------------------------------------------
initial begin reset_n = 0; clock = 0; #3.0 reset_n = 1; #3000 $finish; end
initial begin $dumpfile("tb.vcd"); $dumpvars(0, tb); $readmemh("memory.hex", m, 0); end
// -----------------------------------------------------------------------------
reg  [15:0] m[256*1024];
// -----------------------------------------------------------------------------
wire [19:0] a;
reg  [ 7:0] i;
wire [ 7:0] o;
wire        w;
// -----------------------------------------------------------------------------
always @(negedge clock) begin if (w) m[a] <= o; #0.3 i <= m[a]; end
// -----------------------------------------------------------------------------
c86 T1
(
    .clock      (clock),
    .reset_n    (reset_n),
    .ce         (1'b1),
    .a          (a),
    .i          (i),
    .o          (o),
    .w          (w)
);
// -----------------------------------------------------------------------------
endmodule
