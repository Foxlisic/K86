`timescale 10ns / 1ns
module tb;
// ---------------------------------------------------------------------
reg         clock, clock25, reset_n;
always #0.5 clock       = ~clock;
always #2.0 clock25     = ~clock25;
// ---------------------------------------------------------------------
initial begin reset_n = 0; clock = 0; clock25 = 0; #4.0 reset_n = 1; #2500 $finish; end
initial begin $dumpfile("tb.vcd"); $dumpvars(0, tb); $readmemh("tb.hex", m, 0); end
// ---------------------------------------------------------------------
// Контроллер блочной памяти, до 46Кб, но тут будет 1Мб для совместимости
// ---------------------------------------------------------------------
reg  [ 7:0] m[1024*1024];
wire [19:0] a;
wire [ 7:0] i = m[a];
wire [ 7:0] o;
wire        w;
// ---------------------------------------------------------------------
always @(posedge clock) if (w) m[a] <= o;
// ---------------------------------------------------------------------

micro86 Processor
(
    .clock          (clock25),
    .reset_n        (reset_n),
    .ce             (1'b1),
    .a              (a),
    .i              (i),
    .o              (o),
    .w              (w)
);

endmodule
